module testSerial(output tx, input rx);
  assign tx = rx;
endmodule